// This file is a dummy module for simulation when a pad frame
//   including instantiated corners is used
module PCORNER () ;
endmodule
